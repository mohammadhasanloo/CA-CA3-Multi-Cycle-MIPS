module Memory (input clk,input [31:0] Address, Write_data , input Mem_read , Mem_write , output reg [31:0] Mem_read_value) ;
	reg [31:0] Mem_data [0:4095];
	// Read Data Memory

	initial $readmemb("memory.mem",Mem_data);

	// For Testbench
	wire [31:0] max_element;
	wire [31:0] max_element_i;
	assign max_element_memory = Mem_data[2000];
	assign max_element_i_memory = Mem_data[2004];

	always @(posedge clk) begin
		if( Mem_write )
			Mem_data[Address] <= Write_data;
	end

	assign Mem_read_value = (Mem_read) ? Mem_data[Address] : Mem_read_value;

endmodule